`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: California State University,Chico
// Engineer: Yolanda Reyes #011234614
// 
// Create Date: 02/28/2025 08:23:10 PM
// Design Name: 32-bit Division ALU module with ready bit and clock
// Module Name: divALU32
// Project Name: Homework 0
// Target Devices: That one Basys thing
// Tool Versions: After all this time still a good question...
// Description: Homework 0 purpose is to perform timing and slack analysis
// 
// Dependencies: Electricity, generated from combusting long dead conifers and dinosaurs 
//               or if we are lucky provided by Ehecatl and/or Xiuhcoatl
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module divALU32(                        // Module for performing 32-bit division
    input logic clk,                    // Clock Input
    input logic reset,                  // Enables system to initialize to a known state!
    input logic dividend_in [31:0],     // The value that gets divided "the top part"
    input logic divisor_in [31:0],      // The value that does the dividing "the bottom part"
    output logic quotient_out [31:0],   // The value that results from the division
    output logic remainder_out [31:0],  // The value that is left over after the division
    output logic ready                  // Ready bit is used to determine if all 32 bits have been computed  
);
                                // Internal registers ensure input and outputs are captured properly
    logic [31:0] dividend;      // Internal values, read only stored in REG dividend    
    logic [31:0] divisor;       // Internal values, read only stored in REG divisor
    logic [31:0] quotient;      // Internal values, read only stored in REG quotient
    logic [31:0] remainder;     // Internal values, read only stored in REG remainder
    logic [5:0]  count;         // Internal value, read only to set ready bit @ 33rd iteration
    logic [31:0] temp;          // For temperary values generated by operations
    
    typedef enum logic [2:0]{   // Using enumeration type for state machina implementation
        RESET,                  // State that initializes to known values, all REGs = 0
        SUBTRACT,               // State that performs initial subtraction: Remainder = Remainder - Divisor
        QSHIFT,                 // State that performs the shifting of the quotient REG and sets LSB! Remainder <0 ? LSB =1 : LSB=0
        DSHIFT,                 // State that performs the right by 1-bit shifting of the divisor REG! 
        DONE                    // State that sets the ready bit, do we transition to a reset state?
    }stateMachina_t;
    stateMachina_t current_state, next_state;         // Global module variables associated with stateMachina 
    
    always_ff@(posedge clk or posedge reset) begin  // Flip-Flop to deploy stateMachina for ALU division
        if(reset)begin                              // Reset state ensures initialization with known values executes
            dividend  <= 32'b00000000;              // Set all the internal 32-bit REGs == 0
            divisor   <= 32'b00000000;
            quotient  <= 32'b00000000;
            remainder <= 32'b00000000;
        end else begin                              // This line executes if stateMachina is NOT in reset mode
            current_state = next_state;             // Set the current state to the next state at the positive edge of the clock
        end
        
        case(state)               // Case statements evaluate what the current state is and then execute related codes
           SUBTRACT: begin        // Subtract the divisor REG from the Remainder REG and save the result in Remainder REG
                remainder =  remainder - divisor;
                count++;          // Accumulate how many bits computed so far
                next_state = QSHIFT;    // The next state will be evaluated on the next positive edge of the clock cycle
           end
           
           QSHIFT: begin          // Remainder < 0 ? LSB == 0 : LSB == 1 
                if(remainder < 0) begin     
                    remainder  <=  divisor + remainder;
                    quotient   <= (quotient << 1);    // Shifting to the left 1 bit will pad LSB w/0!
                    count++;                          // Accumulate how many bits computed so far
                    next_state <= DSHIFT;             // The next state will be evaluated on the next positive edge of the clock cycle
                end else begin                        // Shifting to the left 1 bit will pad LSB w/0, the | 1 operation...
                    quotient   <= (quotient << 1) | 1;// Will pad the LSB w/1 since 0 + 1 = 1!
                    count++;                          // Accumulate how many bits computed so far
                    next_state <= DSHIFT;             // The next state will be evaluated on the next positive edge of the clock cycle
                end
           end
           
           DSHIFT: begin                    // Divisor shift 
                divisor = (divisor >> 1);   // Shift the divisor to the right 1-bit
                count++;                    // Accumulate how many bits computed so far
                next_state <= (count == 32) ? DONE : SUBTRACT;  // The next state will be evaluated on the next positive edge of the clock cycle
           end
           
           DONE: begin          // Set the ready bit to signal the ALU has completed computation of the 32-bit division
                ready = 1; 
                next_state <= RESET;    // Will this execute correctly?     
           end 
        endcase
    
endmodule
